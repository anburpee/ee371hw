/* Testbench for Homework 1 Problem 1 */
module hw1p1_tb();

	// for you to implement

	initial begin
	
		// for you to implement
		
	end  // initial
	
endmodule  // hw1p1_tb
