/* Testbench for Homework 1 Problem 2 */
module hw1p2_tb();

	// for you to implement

	initial begin
	
		// for you to implement
		
	end  // initial
	
endmodule  // hw1p2_tb
